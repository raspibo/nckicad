* EESchema Netlist Version 1.1 (Spice format) creation date: mer 29 apr 2015 19:02:55 CEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
IC1  Net-_IC1-Pad1_ Net-_IC1-Pad2_ Net-_IC1-Pad3_ GND GND Net-_IC1-Pad6_ Net-_IC1-Pad7_ VCC Net-_IC1-Pad9_ Net-_IC1-Pad10_ Net-_IC1-Pad11_ GND GND Net-_IC1-Pad14_ Net-_IC1-Pad15_ +5V L293D		
P3  Net-_IC1-Pad6_ Net-_IC1-Pad3_ CONN_01X02		
P4  Net-_IC1-Pad9_ MOTOR2_ENABLE		
P2  Net-_IC1-Pad1_ MOTOR1_ENABLE		
Q1  Net-_Q1-Pad1_ Net-_IC1-Pad7_ GND Q_NPN_BCE		
R2  +5V Net-_IC1-Pad7_ R		
R1  Net-_IC1-Pad2_ Net-_Q1-Pad1_ R		
P1  Net-_IC1-Pad2_ MOTOR1_DIRECTION		
P5  Net-_IC1-Pad11_ Net-_IC1-Pad14_ CONN_01X02		
Q2  Net-_Q2-Pad1_ Net-_IC1-Pad10_ GND Q_NPN_BCE		
R3  +5V Net-_IC1-Pad10_ R		
R4  Net-_IC1-Pad15_ Net-_Q2-Pad1_ R		
P6  Net-_IC1-Pad15_ MOTOR2_DIRECTION		
P8  +5V CONN_01X01		
P7  VCC CONN_01X01		
P9  GND CONN_01X01		

.end
